magic
tech sky130A
magscale 1 2
timestamp 1707327043
<< viali >>
rect 1128 2926 1272 3046
rect 1676 1846 1826 1978
<< metal1 >>
rect 100 3204 2904 3402
rect 732 3190 932 3204
rect 1098 3046 1300 3204
rect 1098 2926 1128 3046
rect 1272 2926 1300 3046
rect 1098 2814 1300 2926
rect 638 2718 880 2734
rect 638 2636 684 2718
rect 846 2636 880 2718
rect 638 2606 880 2636
rect 378 2466 578 2482
rect -138 2444 1120 2466
rect -138 2350 -92 2444
rect 16 2350 386 2444
rect -138 2328 386 2350
rect 542 2442 1120 2444
rect 542 2350 1028 2442
rect 1112 2350 1120 2442
rect 542 2328 1120 2350
rect 378 2282 578 2328
rect 1506 2100 1574 2106
rect 664 2062 864 2090
rect 664 1926 690 2062
rect 840 1926 864 2062
rect 1506 2048 1508 2100
rect 1572 2048 1574 2100
rect 1506 2040 1574 2048
rect 664 1890 864 1926
rect 1394 1972 1490 1994
rect 1394 1868 1418 1972
rect 1394 1850 1490 1868
rect 1596 1978 2202 2000
rect 1596 1846 1676 1978
rect 1826 1846 2202 1978
rect 1596 1830 2202 1846
rect 640 1396 840 1406
rect 2000 1396 2198 1830
rect -4 1198 2800 1396
<< via1 >>
rect 684 2636 846 2718
rect -92 2350 16 2444
rect 386 2328 542 2444
rect 1028 2350 1112 2442
rect 690 1926 840 2062
rect 1508 2048 1572 2100
rect 1418 1868 1490 1972
<< metal2 >>
rect -98 2736 452 2792
rect -96 2444 40 2736
rect 632 2718 892 2744
rect 632 2636 684 2718
rect 846 2636 892 2718
rect -96 2350 -92 2444
rect 16 2350 40 2444
rect -96 2328 40 2350
rect 378 2444 578 2482
rect 378 2328 386 2444
rect 542 2328 578 2444
rect 378 2282 578 2328
rect 632 2062 892 2636
rect 1020 2442 1690 2466
rect 1020 2350 1028 2442
rect 1112 2350 1690 2442
rect 1020 2326 1690 2350
rect 632 1926 690 2062
rect 840 2000 892 2062
rect 1506 2100 1574 2326
rect 1506 2048 1508 2100
rect 1572 2048 1574 2100
rect 1506 2040 1574 2048
rect 840 1972 1490 2000
rect 840 1926 1418 1972
rect 632 1868 1418 1926
rect 632 1838 1490 1868
use sky130_fd_pr__pfet_01v8_XPMKZ5  XM1
timestamp 1707214941
transform 0 1 1491 -1 0 2764
box -246 -1219 246 1219
use sky130_fd_pr__nfet_01v8_PVEW3M  XM2
timestamp 1707214941
transform 1 0 1540 0 1 1918
box -246 -310 246 310
<< labels >>
flabel metal1 378 2282 578 2482 0 FreeSans 256 0 0 0 Vin
port 0 nsew
flabel metal1 640 1206 840 1406 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 732 3190 932 3390 0 FreeSans 256 0 0 0 VDD
port 2 nsew
flabel metal1 664 1890 864 2090 0 FreeSans 256 0 0 0 Vout
port 3 nsew
<< end >>
